package common is 

    type int_vector is array (0 to 3) of integer;
    type states_t is (HOLA, NUM1, NUM2, CHECK, BIEN, ERROR, PR1, PR2);

end common;

package body common is
end common;